module datapath
#(
    parameter WORD_SIZE = 32
)
(
    input wire clock
);
    
    // IMPORT DATA_PATH TEST AND SET IT AS A PROPER DATAPATH MODULE

endmodule